module vga_pic(
input wire vga_clk , //输入工作时钟,频率25MHz
input wire sys_rst_n , //输入复位信号,低电平有效
input wire [9:0] pix_x , //输入有效显示区域像素点X轴坐标
input wire [9:0] pix_y , //输入有效显示区域像素点Y轴坐标

output reg [15:0] pix_data //输出像素点色彩信息

);

////
//\* Parameter and Internal Signal \//
////
//parameter define
parameter CHAR_B_H= 10'd192 , //字符开始X轴坐标
CHAR_B_V= 10'd208 ; //字符开始Y轴坐标

parameter CHAR_W = 10'd256 , //字符宽度
CHAR_H = 10'd64 ; //字符高度

parameter BLACK = 16'h0000, //黑色
WHITE = 16'hFFFF, //白色
GOLDEN = 16'hFEC0; //金色

//wire define
wire [9:0] char_x ; //字符显示X轴坐标
wire [9:0] char_y ; //字符显示Y轴坐标

//reg define
reg [255:0] char [63:0] ; //字符数据

////
//\* Main Code \//
////

//字符显示坐标
assign char_x = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
? (pix_x - CHAR_B_H) : 10'h3FF;
assign char_y = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
? (pix_y - CHAR_B_V) : 10'h3FF;

//char:字符数据
always@(posedge vga_clk)
begin
char[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[3] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[4] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[5] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[6] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[7] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[8] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[9] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[10] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[11] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[12] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[13] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[14] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[15] <= 256'h000000000000000000000000000000000000007FF80000000000000000000000;
char[16] <= 256'h00000000001FFF80001FFF801FFC000FFC0003FFFFC00FFFFFFFFFC000000000;
char[17] <= 256'h00000000001FFF80001FFF801FFC000FFC000FFFFFF80FFFFFFFFFC000000000;
char[18] <= 256'h00000000001FFFC0003FFF801FFC000FFC001FFFFFF80FFFFFFFFFC000000000;
char[19] <= 256'h00000000001FFFC0003FFF801FFC000FFC003FFFFFF80FFFFFFFFFC000000000;
char[20] <= 256'h00000000001FFFC0007FFF801FFC000FFC007FFFFFF80FFFFFFFFFC000000000;
char[21] <= 256'h00000000001FFFE0007FFF801FFC000FFC00FFFFFFF80FFFFFFFFFC000000000;
char[22] <= 256'h00000000001FFFE000FFFF801FFC000FFC00FFFFFFF80FFFFFFFFFC000000000;
char[23] <= 256'h00000000001FFFF000FFFF801FFC000FFC00FFF007F80FFFFFFFFFC000000000;
char[24] <= 256'h00000000001FFFF000FFFF801FFC000FFC01FFC0007800003FF0000000000000;
char[25] <= 256'h00000000001FFFF801FFFF801FFC000FFC01FF80001000003FF0000000000000;
char[26] <= 256'h00000000001FFFF801FFFF801FFC000FFC01FF80000000003FF0000000000000;
char[27] <= 256'h00000000001FFFF803FFFF801FFC000FFC01FF80000000003FF0000000000000;
char[28] <= 256'h00000000001FFBFC03FDFF801FFC000FFC01FF80000000003FF0000000000000;
char[29] <= 256'h00000000001FFBFC07FDFF801FFC000FFC01FF80000000003FF0000000000000;
char[30] <= 256'h00000000001FF9FE07F9FF801FFC000FFC01FFE0000000003FF0000000000000;
char[31] <= 256'h00000000001FF9FE07F9FF801FFC000FFC00FFFE000000003FF0000000000000;
char[32] <= 256'h00000000001FF9FF0FF1FF801FFC000FFC00FFFFF00000003FF0000000000000;
char[33] <= 256'h00000000001FF8FF0FF1FF801FFC000FFC00FFFFFE0000003FF0000000000000;
char[34] <= 256'h00000000001FF8FF1FE1FF801FFC000FFC007FFFFF8000003FF0000000000000;
char[35] <= 256'h00000000001FF87F9FE1FF801FFC000FFC003FFFFFE000003FF0000000000000;
char[36] <= 256'h00000000001FF87FBFE1FF801FFC000FFC001FFFFFF000003FF0000000000000;
char[37] <= 256'h00000000001FF83FFFC1FF801FFC000FFC000FFFFFF800003FF0000000000000;
char[38] <= 256'h00000000001FF83FFFC1FF801FFC000FFC0003FFFFFC00003FF0000000000000;
char[39] <= 256'h00000000001FF83FFF81FF801FFC000FFC00007FFFFC00003FF0000000000000;
char[40] <= 256'h00000000001FF81FFF81FF801FFC000FFC000007FFFE00003FF0000000000000;
char[41] <= 256'h00000000001FF81FFF01FF801FFC000FFC0000007FFE00003FF0000000000000;
char[42] <= 256'h00000000001FF80FFF01FF801FFC000FFC0000001FFE00003FF0000000000000;
char[43] <= 256'h00000000001FF80FFF01FF801FFC000FFC0000000FFE00003FF0000000000000;
char[44] <= 256'h00000000001FF807FE01FF801FFC001FFC00000007FE00003FF0000000000000;
char[45] <= 256'h00000000001FF807FE01FF800FFC001FFC00000007FE00003FF0000000000000;
char[46] <= 256'h00000000001FF807FC01FF800FFE001FFC01000007FE00003FF0000000000000;
char[47] <= 256'h00000000001FF803FC01FF800FFE003FF801E00007FE00003FF0000000000000;
char[48] <= 256'h00000000001FF803F801FF800FFF007FF801F8000FFE00003FF0000000000000;
char[49] <= 256'h00000000001FF8000001FF8007FFC0FFF801FF803FFC00003FF0000000000000;
char[50] <= 256'h00000000001FF8000001FF8007FFFFFFF001FFFFFFFC00003FF0000000000000;
char[51] <= 256'h00000000001FF8000001FF8003FFFFFFF001FFFFFFFC00003FF0000000000000;
char[52] <= 256'h00000000001FF8000001FF8003FFFFFFE001FFFFFFF800003FF0000000000000;
char[53] <= 256'h00000000001FF8000001FF8001FFFFFFC001FFFFFFF000003FF0000000000000;
char[54] <= 256'h00000000001FF8000001FF8000FFFFFF8001FFFFFFE000003FF0000000000000;
char[55] <= 256'h00000000001FF8000001FF80003FFFFF00007FFFFFC000003FF0000000000000;
char[56] <= 256'h00000000001FF8000001FF80000FFFFC00000FFFFF0000003FF0000000000000;
char[57] <= 256'h0000000000000000000000000001FFC00000007FF80000000000000000000000;
char[58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
end

 //pix_data:输出像素点色彩信息,根据当前像素点坐标指定当前像素点颜色数据
 always@(posedge vga_clk or negedge sys_rst_n)
 if(sys_rst_n == 1'b0)
 pix_data <= BLACK;
 else if((((pix_x >= (CHAR_B_H - 1'b1))
 && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
 && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
 && (char[char_y][10'd255 - char_x] == 1'b1))
 pix_data <= GOLDEN;
 else
 pix_data <= BLACK;

 endmodule